module main();
initial
  begin
    $hello;
    $display("Hi there");
    $finish;
  end

endmodule
